module full_add ( 
    input a, b, cin,
    output sum, cout );

    // write code here


endmodule