module lut_top (
<<<<<<< HEAD
    input clk,
    input enable,
    input S,
    input A, B, C,
    output Z 
);
    
    reg [7:0] Q;
    
    assign Z = Q[{A, B, C}];
   	
    always @(posedge clk) begin
        
        if (enable) Q <= {Q[6:0], S};
       
    end
=======

);
    

>>>>>>> 0903dde (review 3 labs)
endmodule
