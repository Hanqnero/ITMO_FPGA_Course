module full_add ( 
    input a, b, cin,
    output sum, cout );

<<<<<<< HEAD
    assign sum = a != b != cin;
    assign cout = a && b || a && cin || b && cin;
=======
    // write code here
>>>>>>> 0903dde (review 3 labs)

endmodule