module Analyse (
    input a, b, c, d,
    output q
);
    assign q = b | c;
endmodule